//lut查找表 256
module lut_256(clk,rst,addr,out);
 input clk;
 input rst;
 input [7:0] addr;
 output[15:0] out;
 
 reg[15:0] out_tmp;
 
always @ ( posedge clk or negedge rst )
        if(!rst)
           out_tmp <= 16'd0;
        else
           case(addr)
                
                0,1  :   out_tmp <= 16'd0;
                2    :   out_tmp <= 16'd1;
                3    :   out_tmp <= 16'd2;
                4    :   out_tmp <= 16'd4;
                5    :   out_tmp <= 16'd6;
                6    :   out_tmp <= 16'd9;
                7    :   out_tmp <= 16'd12;
                8    :   out_tmp <= 16'd16;
                9    :   out_tmp <= 16'd20;
                10   :   out_tmp <= 16'd25;
                11   :   out_tmp <= 16'd30;
                12   :   out_tmp <= 16'd36;
                13   :   out_tmp <= 16'd42;
                14   :   out_tmp <= 16'd49;
                15   :   out_tmp <= 16'd56;
                16   :   out_tmp <= 16'd64;
                17   :   out_tmp <= 16'd72;
                18   :   out_tmp <= 16'd81;
                19   :   out_tmp <= 16'd90;
                20   :   out_tmp <= 16'd100;
                21   :   out_tmp <= 16'd110;
                22   :   out_tmp <= 16'd121;
                23   :   out_tmp <= 16'd132;
                24   :   out_tmp <= 16'd144;
                25   :   out_tmp <= 16'd156;
                26   :   out_tmp <= 16'd169;
                27   :   out_tmp <= 16'd182;
                28   :   out_tmp <= 16'd196;
                29   :   out_tmp <= 16'd210;
                30   :   out_tmp <= 16'd225;
                31   :   out_tmp <= 16'd240;
                32   :   out_tmp <= 16'd256;
                33   :   out_tmp <= 16'd272;
                34   :   out_tmp <= 16'd289;
                35   :   out_tmp <= 16'd306;
                36   :   out_tmp <= 16'd324;
                37   :   out_tmp <= 16'd342;
                38   :   out_tmp <= 16'd361;
                39   :   out_tmp <= 16'd380;
                40   :   out_tmp <= 16'd400;
                41   :   out_tmp <= 16'd420;
                42   :   out_tmp <= 16'd441;
                43   :   out_tmp <= 16'd462;
                44   :   out_tmp <= 16'd484;
                45   :   out_tmp <= 16'd506;
                46   :   out_tmp <= 16'd529;
                47   :   out_tmp <= 16'd552;
                48   :   out_tmp <= 16'd576;
                49   :   out_tmp <= 16'd600;
                50   :   out_tmp <= 16'd625;
                51   :   out_tmp <= 16'd650;
                52   :   out_tmp <= 16'd676;
                53   :   out_tmp <= 16'd702;
                54   :   out_tmp <= 16'd729;
                55   :   out_tmp <= 16'd756;
                56   :   out_tmp <= 16'd784;
                57   :   out_tmp <= 16'd812;
                58   :   out_tmp <= 16'd841;
                59   :   out_tmp <= 16'd870;
                60   :   out_tmp <= 16'd900;
                61   :   out_tmp <= 16'd930;
                62   :   out_tmp <= 16'd961;
                63   :   out_tmp <= 16'd992;
                64   :   out_tmp <= 16'd1024;
                65   :   out_tmp <= 16'd1056;
                66   :   out_tmp <= 16'd1089;
                67   :   out_tmp <= 16'd1122;
                68   :   out_tmp <= 16'd1156;
                69   :   out_tmp <= 16'd1190;
                70   :   out_tmp <= 16'd1225;
                71   :   out_tmp <= 16'd1260;
                72   :   out_tmp <= 16'd1296;
                73   :   out_tmp <= 16'd1332;
                74   :   out_tmp <= 16'd1369;
                75   :   out_tmp <= 16'd1406;
                76   :   out_tmp <= 16'd1444;
                77   :   out_tmp <= 16'd1482;
                78   :   out_tmp <= 16'd1521;
                79   :   out_tmp <= 16'd1560;
                80   :   out_tmp <= 16'd1600;
                81   :   out_tmp <= 16'd1640;
                82   :   out_tmp <= 16'd1681;
                83   :   out_tmp <= 16'd1722;
                84   :   out_tmp <= 16'd1764;
                85   :   out_tmp <= 16'd1806;
                86   :   out_tmp <= 16'd1849;
                87   :   out_tmp <= 16'd1892;
                88   :   out_tmp <= 16'd1936;
                89   :   out_tmp <= 16'd1980;
                90   :   out_tmp <= 16'd2025;
                91   :   out_tmp <= 16'd2070;
                92   :   out_tmp <= 16'd2116;
                93   :   out_tmp <= 16'd2162;
                94   :   out_tmp <= 16'd2209;
                95   :   out_tmp <= 16'd2256;
                96   :   out_tmp <= 16'd2304;
                97   :   out_tmp <= 16'd2352;
                98   :   out_tmp <= 16'd2401;
                99   :   out_tmp <= 16'd2450;
                100  :   out_tmp <= 16'd2500;
                101  :   out_tmp <= 16'd2550;
                102  :   out_tmp <= 16'd2601;
                103  :   out_tmp <= 16'd2652;
                104  :   out_tmp <= 16'd2704;
                105  :   out_tmp <= 16'd2756;
                106  :   out_tmp <= 16'd2809;
                107  :   out_tmp <= 16'd2862;
                108  :   out_tmp <= 16'd2916;
                109  :   out_tmp <= 16'd2970;
                110  :   out_tmp <= 16'd3025;
                111  :   out_tmp <= 16'd3080;
                112  :   out_tmp <= 16'd3136;
                113  :   out_tmp <= 16'd3192;
                114  :   out_tmp <= 16'd3249;
                115  :   out_tmp <= 16'd3306;
                116  :   out_tmp <= 16'd3364;
                117  :   out_tmp <= 16'd3422;
                118  :   out_tmp <= 16'd3481;
                119  :   out_tmp <= 16'd3540;
                120  :   out_tmp <= 16'd3600;
                121  :   out_tmp <= 16'd3660;
                122  :   out_tmp <= 16'd3721;
                123  :   out_tmp <= 16'd3782;
                124  :   out_tmp <= 16'd3844;
                125  :   out_tmp <= 16'd3906;
                126  :   out_tmp <= 16'd3969;
                127  :   out_tmp <= 16'd4032;
                128  :   out_tmp <= 16'd4096;
                129  :   out_tmp <= 16'd4160;
                130  :   out_tmp <= 16'd4225;
                131  :   out_tmp <= 16'd4290;
                132  :   out_tmp <= 16'd4356;
                133  :   out_tmp <= 16'd4422;
                134  :   out_tmp <= 16'd4489;
                135  :   out_tmp <= 16'd4556;
                136  :   out_tmp <= 16'd4624;
                137  :   out_tmp <= 16'd4692;
                138  :   out_tmp <= 16'd4761;
                139  :   out_tmp <= 16'd4830;
                140  :   out_tmp <= 16'd4900;
                141  :   out_tmp <= 16'd4970;
                142  :   out_tmp <= 16'd5041;
                143  :   out_tmp <= 16'd5112;
                144  :   out_tmp <= 16'd5184;
                145  :   out_tmp <= 16'd5256;
                146  :   out_tmp <= 16'd5329;
                147  :   out_tmp <= 16'd5402;
                148  :   out_tmp <= 16'd5476;
                149  :   out_tmp <= 16'd5550;
                150  :   out_tmp <= 16'd5625;
                151  :   out_tmp <= 16'd5700;
                152  :   out_tmp <= 16'd5776;
                153  :   out_tmp <= 16'd5852;
                154  :   out_tmp <= 16'd5929;
                155  :   out_tmp <= 16'd6006;
                156  :   out_tmp <= 16'd6084;
                157  :   out_tmp <= 16'd6162;
                158  :   out_tmp <= 16'd6241;
                159  :   out_tmp <= 16'd6320;
                160  :   out_tmp <= 16'd6400;
                161  :   out_tmp <= 16'd6480;
                162  :   out_tmp <= 16'd6561;
                163  :   out_tmp <= 16'd6642;
                164  :   out_tmp <= 16'd6724;
                165  :   out_tmp <= 16'd6806;
                166  :   out_tmp <= 16'd6889;
                167  :   out_tmp <= 16'd6972;
                168  :   out_tmp <= 16'd7056;
                169  :   out_tmp <= 16'd7140;
                170  :   out_tmp <= 16'd7225;
                171  :   out_tmp <= 16'd7310;
                172  :   out_tmp <= 16'd7396;
                173  :   out_tmp <= 16'd7482;
                174  :   out_tmp <= 16'd7569;
                175  :   out_tmp <= 16'd7656;
                176  :   out_tmp <= 16'd7744;
                177  :   out_tmp <= 16'd7832;
                178  :   out_tmp <= 16'd7921;
                179  :   out_tmp <= 16'd8010;
                180  :   out_tmp <= 16'd8100;
                181  :   out_tmp <= 16'd8190;
                182  :   out_tmp <= 16'd8281;
                183  :   out_tmp <= 16'd8372;
                184  :   out_tmp <= 16'd8464;
                185  :   out_tmp <= 16'd8556;
                186  :   out_tmp <= 16'd8649;
                187  :   out_tmp <= 16'd8742;
                188  :   out_tmp <= 16'd8836;
                189  :   out_tmp <= 16'd8930;
                190  :   out_tmp <= 16'd9025;
                191  :   out_tmp <= 16'd9120;
                192  :   out_tmp <= 16'd9216;
                193  :   out_tmp <= 16'd9312;
                194  :   out_tmp <= 16'd9409;
                195  :   out_tmp <= 16'd9506;
                196  :   out_tmp <= 16'd9604;
                197  :   out_tmp <= 16'd9702;
                198  :   out_tmp <= 16'd9801;
                199  :   out_tmp <= 16'd9900;
                200  :   out_tmp <= 16'd10000;
                201  :   out_tmp <= 16'd10100;
                202  :   out_tmp <= 16'd10201;
                203  :   out_tmp <= 16'd10302;
                204  :   out_tmp <= 16'd10404;
                205  :   out_tmp <= 16'd10506;
                206  :   out_tmp <= 16'd10609;
                207  :   out_tmp <= 16'd10712;
                208  :   out_tmp <= 16'd10816;
                209  :   out_tmp <= 16'd10920;
                210  :   out_tmp <= 16'd11025;
                211  :   out_tmp <= 16'd11130;
                212  :   out_tmp <= 16'd11236;
                213  :   out_tmp <= 16'd11342;
                214  :   out_tmp <= 16'd11449;
                215  :   out_tmp <= 16'd11556;
                216  :   out_tmp <= 16'd11664;
                217  :   out_tmp <= 16'd11772;
                218  :   out_tmp <= 16'd11881;
                219  :   out_tmp <= 16'd11990;
                220  :   out_tmp <= 16'd12100;
                221  :   out_tmp <= 16'd12210;
                222  :   out_tmp <= 16'd12321;
                223  :   out_tmp <= 16'd12432;
                224  :   out_tmp <= 16'd12544;
                225  :   out_tmp <= 16'd12656;
                226  :   out_tmp <= 16'd12769;
                227  :   out_tmp <= 16'd12882;
                228  :   out_tmp <= 16'd12996;
                229  :   out_tmp <= 16'd13100;
                230  :   out_tmp <= 16'd13225;
                231  :   out_tmp <= 16'd13340;
                232  :   out_tmp <= 16'd13456;
                233  :   out_tmp <= 16'd13572;
                234  :   out_tmp <= 16'd13689;
                235  :   out_tmp <= 16'd13806;
                236  :   out_tmp <= 16'd13924;
                237  :   out_tmp <= 16'd14042;
                238  :   out_tmp <= 16'd14161;
                239  :   out_tmp <= 16'd14280;
                240  :   out_tmp <= 16'd14400;
                241  :   out_tmp <= 16'd14520;
                242  :   out_tmp <= 16'd14641;
                243  :   out_tmp <= 16'd14762;
                244  :   out_tmp <= 16'd14884;
                245  :   out_tmp <= 16'd15006;
                246  :   out_tmp <= 16'd15129;
                247  :   out_tmp <= 16'd15252;
                248  :   out_tmp <= 16'd15376;
                249  :   out_tmp <= 16'd15500;
                250  :   out_tmp <= 16'd15625;
                251  :   out_tmp <= 16'd15750;
                252  :   out_tmp <= 16'd15876;
                253  :   out_tmp <= 16'd16002;
                254  :   out_tmp <= 16'd16129;
                255  :   out_tmp <= 16'd16256;
        
        endcase
assign out=out_tmp;
endmodule